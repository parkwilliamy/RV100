`timescale 1ns/1ps

module StallUnit (
    input EX_MemRead,
    input [4:0] EX_rd, ID_rs1, ID_rs2,
    input [2:0] ID_ValidReg,
    output reg Stall
);

    always @ (*) begin

        if (EX_MemRead) begin

            Stall = (((EX_rd == ID_rs1) && ID_ValidReg[1])) || ((EX_rd == ID_rs2) && ID_ValidReg[2]);

        end

        else Stall = 0;

    end


endmodule